RL Load SCR circuit
