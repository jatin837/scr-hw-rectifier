RL load SCR
.include include/thy.sub
