RL load SCR
